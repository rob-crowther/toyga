Untitled

R0 n2 0 820000
C1 n3 0 3.9e-11
R1 n3 n1 51000000
R2 n1 n4 220000
R3 0 n4 6200000
R4 n4 n3 13000
L1 n6 0 1.3e-08
C2 n3 n4 3.9e-07

VIN n1 0 DC 5 AC 1 PULSE(0 1 0.0000005 0.000000000001 0.000000000001 1 2) 

.op
.ac lin 1000 100000 100
.plot ac vdb(n1) xlog
.end
